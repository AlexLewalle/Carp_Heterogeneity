-85.8318            # Vm
1                   # Lambda
0                   # delLambda
2.9142e-06          # Tension
-                   # K_e
-                   # Na_e
-                   # Ca_e
7.97028e-05         # Iion
-                   # tension_component
TT2_Cai
2.38899             # CaSR
0.000193312         # CaSS
0.0823333           # Ca_i
3.11213e-05         # D
0.976267            # F
0.999293            # F2
0.999747            # FCaSS
3.98e-05            # GCaL
0.153               # Gkr
0.392               # Gks
0.294               # Gto
0.76102             # H
0.760739            # J
138.087             # K_i
0.00150933          # M
7.57291             # Na_i
2.18602e-08         # R
0.989506            # R_
0.999973            # S
0.000194378         # Xr1
0.477427            # Xr2
0.00313223          # Xs

LandStress
0                   # Q_1
0                   # Q_2
0.0104987           # TRPN
2.42848e-08         # xb
0                   # __Ca_i_local

