-85.4192            # Vm
1                   # Lambda
0                   # delLambda
2.21177e-05         # Tension
-                   # K_e
-                   # Na_e
-                   # Ca_e
9.58674e-05         # Iion
-                   # tension_component
TT2_Cai
3.35309             # CaSR
0.000210233         # CaSS
0.101105            # Ca_i
3.28817e-05         # D
0.976433            # F
0.999264            # F2
0.999745            # FCaSS
3.98e-05            # GCaL
0.153               # Gkr
0.392               # Gks
0.294               # Gto
0.75005             # H
0.749607            # J
136.267             # K_i
0.00164781          # M
8.68579             # Na_i
2.34171e-08         # R
0.989115            # R_
0.999973            # S
0.000206442         # Xr1
0.473141            # Xr2
0.00322439          # Xs

LandStress
0                   # Q_1
0                   # Q_2
0.0157463           # TRPN
1.84313e-07         # xb
0                   # __Ca_i_local

