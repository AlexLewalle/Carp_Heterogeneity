84.395              # Vm
1                   # Lambda
0                   # delLambda
119.373             # Tension
-                   # K_e
-                   # Na_e
-                   # Ca_e
0.0112987           # Iion
-                   # tension_component
TT2_Cai
2.34796             # CaSR
1.09946             # CaSS
1000                # Ca_i
0.999997            # D
0.0105963           # F
0.330046            # F2
0.401242            # FCaSS
3.98e-05            # GCaL
0.153               # Gkr
0.392               # Gks
0.294               # Gto
5.87954e-19         # H
5.8823e-19          # J
131.75              # K_i
1                   # M
28.0395             # Na_i
0.999981            # R
0.0657902           # R_
8.50041e-10         # S
1                   # Xr1
0.000758441         # Xr2
0.99815             # Xs

LandHumanStress
0.999999            # TRPN
0.00522476          # TmBlocked
0.248694            # XS
0.373041            # XW
0                   # ZETAS
0                   # ZETAW
0                   # __Ca_i_local

