-4.0772             # Vm
1                   # Lambda
0                   # delLambda
5.78575e-07         # Tension
-                   # K_e
-                   # Na_e
-                   # Ca_e
0.512746            # Iion
-                   # tension_component
TT2_Cai
1.27809             # CaSR
0.018539            # CaSS
0.07                # Ca_i
0.643082            # D
0.207106            # F
0.332921            # F2
0.889367            # FCaSS
3.98e-05            # GCaL
0.153               # Gkr
0.392               # Gks
0.294               # Gto
1.24891e-08         # H
1.00934e-08         # J
138.267             # K_i
0.994258            # M
7.64274             # Na_i
0.0274656           # R
0.744082            # R_
0.0228908           # S
0.994347            # Xr1
0.0277576           # Xr2
0.194534            # Xs

LandStress
0                   # Q_1
0                   # Q_2
0.00759808          # TRPN
4.82146e-09         # xb
0                   # __Ca_i_local

