-85.1192            # Vm
1                   # Lambda
0                   # delLambda
0.0110933           # Tension
-                   # K_e
-                   # Na_e
-                   # Ca_e
0.00302465          # Iion
0                   # tension_component
TT2_Cai_init
0.13553             # Ca_i
3.90357             # CaSR
0.000390854         # CaSS
0.904553            # R_
2.8959e-07          # O
7.96934             # Na_i
137.474             # K_i
0.00176341          # M
0.740048            # H
0.668894            # J
0.0173138           # Xr1
0.469827            # Xr2
0.0147276           # Xs
2.47707e-08         # R
0.999995            # S
3.43115e-05         # D
0.72632             # F
0.958372            # F2
0.995453            # FCaSS

LandStress
0                   # Q_1
0                   # Q_2
0.0205164           # TRPN
7.79904e-05         # xb
0                   # __Ca_i_local

