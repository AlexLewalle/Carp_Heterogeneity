-86.0787            # Vm
1                   # Lambda
0                   # delLambda
2.0018e-07          # Tension
-                   # K_e
-                   # Na_e
-                   # Ca_e
7.02765e-05         # Iion
-                   # tension_component
TT2_Cai
1.44171             # CaSR
0.000178208         # CaSS
0.0628352           # Ca_i
3.01135e-05         # D
0.976956            # F
0.999309            # F2
0.999748            # FCaSS
3.98e-05            # GCaL
0.153               # Gkr
0.392               # Gks
0.294               # Gto
0.767411            # H
0.767221            # J
138.277             # K_i
0.00143201          # M
7.64991             # Na_i
2.09788e-08         # R
0.989807            # R_
0.999973            # S
0.000187545         # Xr1
0.479995            # Xr2
0.00307781          # Xs

LandStress
0                   # Q_1
0                   # Q_2
0.00614489          # TRPN
1.66815e-09         # xb
0                   # __Ca_i_local

