-81.6453            # Vm
1                   # Lambda
0                   # delLambda
0.807489            # Tension
-                   # K_e
-                   # Na_e
-                   # Ca_e
0.000533058         # Iion
0                   # tension_component
GPB_Land
6.75947e-07         # C1
0.000620798         # C10
0.0205442           # C11
0.198039            # C12
0.00250135          # C13
0.0606538           # C14
0.0188605           # C15
1.35154e-05         # C2
0.000388903         # C3
0.0117104           # C4
0.258254            # C5
6.07298e-05         # C6
0.00312862          # C7
0.0545955           # C8
0.359934            # C9
0.000350703         # CaM
0.103239            # Ca_i
0.512397            # Ca_sr
0.000192956         # Caj
0.000133056         # Casl
1.14611             # Csqnb
120.327             # Ki
0.00258741          # Myoc
0.136892            # Myom
3.59287             # NaBj
0.783843            # NaBsl
9.0493              # Nai
9.04872             # Naj
9.04904             # Nasl
0.00581863          # O1
0                   # Q_1
0                   # Q_2
2.07956e-07         # RyRi
7.16057e-07         # RyRo
0.774948            # RyRr
0.0786257           # SLHj
0.13695             # SLHsl
0.00811755          # SLLj
0.012327            # SLLsl
0.00255317          # SRB
0.0775398           # TRPN
0.122195            # TnCHc
0.00837978          # TnCHm
0.00542779          # TnCL
2.83308e-06         # d
0.993897            # f
0.0350807           # fcaBj
0.0240456           # fcaBsl
0.632363            # h
0.630237            # j
0.0036461           # m
0.00567697          # xb
0.155557            # xkr
0.00422483          # xks
0.000434241         # xtof
0.0004344           # xtos
0.999986            # ytof
0.526964            # ytos

