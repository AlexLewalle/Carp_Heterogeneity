24.7047             # Vm
1                   # Lambda
0                   # delLambda
0.0009224           # Tension
-                   # K_e
-                   # Na_e
-                   # Ca_e
-0.649676           # Iion
-                   # tension_component
TT2_Cai
1.29122             # CaSR
0.168524            # CaSS
0.0883063           # Ca_i
0.987139            # D
0.954777            # F
0.73323             # F2
0.761929            # FCaSS
3.98e-05            # GCaL
0.153               # Gkr
0.392               # Gks
0.294               # Gto
5.77319e-12         # H
1.92365e-10         # J
138.292             # K_i
0.99976             # M
7.67802             # Na_i
0.655275            # R
0.934399            # R_
0.152383            # S
0.354456            # Xr1
0.0338722           # Xr2
0.00791478          # Xs

LandStress
0                   # Q_1
0                   # Q_2
0.0331136           # TRPN
7.66176e-06         # xb
0                   # __Ca_i_local

